`timescale 1ns / 100ps
/*******************************************************************************
*         (c) Copyright 1997,  National Semiconductor Corporation
*                           ALL RIGHTS RESERVED
********************************************************************************
*                   NATIONAL SEMICONDUCTOR CONFIDENTIAL
********************************************************************************
* *$Id: template_hdl.v,v 1.1 1998/07/09 22:49:34 clk Exp $
* *Name: or2_gea0
*===============================================================================
* *History: $Id$
*    Nov, 27 00 | <marcello@enigma>: V1.00 First edit
*===============================================================================
* *Description:
*
* parent:  (Upward hierarchy) If known
* children:  (downward hierarchy)
*
* *endName
********************************************************************************
********************************************************************************
*        1         2         3         4         5         6         7         8
*2345678901234567890123456789012345678901234567890123456789012345678901234567890
*******************************************************************************/

module or2_gea0 (y, a, b);
   output y; // output
   input a; // first input
   input b; // second input
 
  assign y = (a | b);

endmodule // of or2_gea0

