`timescale 100 ps/100 ps
/*******************************************************************************
*         (c) Copyright 1997,  National Semiconductor Corporation
*                           ALL RIGHTS RESERVED
********************************************************************************
*                   NATIONAL SEMICONDUCTOR CONFIDENTIAL
********************************************************************************
* *$Id: template_hdl.v,v 1.1 1998/07/09 22:49:34 clk Exp $
* *Name: inv_gea1
*===============================================================================
* *History: $Id$
*   Mon Oct 16 11:31:06 MET DST 2000 - v1  marcello      Initial Revision
*===============================================================================
* *Description:
*
* parent:  (Upward hierarchy) If known
* children:  (downward hierarchy)
*
* *endName
********************************************************************************
********************************************************************************
*        1         2         3         4         5         6         7         8
*2345678901234567890123456789012345678901234567890123456789012345678901234567890
*******************************************************************************/
 
module inv_gea1 (y,a);
   output y; // inv_gea1's output
   input  a; // inv_gea1's input
   
   assign y = ~a;
    
 
endmodule  //  End of 'module inv_gea1 ()'

